//----------------------------------------------------------------------------
//
//  Пример 3: Буква в зависимости от кнопки
//
//----------------------------------------------------------------------------

//----------------------------------------------------------------------------
//
// Вариант 1. Выводим букву 'Y' на семисегментный индикатор,
// используя операторы непрерывного присваивания для каждого бита
//
//----------------------------------------------------------------------------

module top_1
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    assign pio [7] = 1'b0;  // a
    assign pio [6] = 1'b1;  // b
    assign pio [5] = 1'b1;  // c
    assign pio [4] = 1'b1;  // d
    assign pio [3] = 1'b0;  // e
    assign pio [2] = 1'b1;  // f
    assign pio [1] = 1'b1;  // g

endmodule

    
//----------------------------------------------------------------------------
//
// Вариант 2. Выводим одну букву P. Присваиваем целым битовым вектором.
// используя операторы непрерывного присваивания для каждого бита
//
//----------------------------------------------------------------------------

module top_2
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    assign pio [7:1] = 7'b1100111;  // abcdefg

endmodule

//----------------------------------------------------------------------------
//
// Вариант 3. Выводим Y или P в зависимости от кнопки 0.
//
//----------------------------------------------------------------------------

module top_3
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    assign pio [7:1] = BTN [0] ? 7'b1100111 /* P */ : 7'b0111011 /* Y */ ;

endmodule

//----------------------------------------------------------------------------
//
// Вариант 4. Выводим Y или P в зависимости от кнопки 0. Кнопка 1 переворачивает букву.
// Способ 1. assign и операция '?'
//
//----------------------------------------------------------------------------

module top_4
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    assign pio [7:1]
        = 
        BTN [1] 
            ? (BTN [0]
                ? 7'b0111101     // перевернутое P
                : 7'b1010111 )   // перевернутое Y
            : (BTN [0]
                ? 7'b1100111     // P
                : 7'b0111011 );  // Y

endmodule

//----------------------------------------------------------------------------
//
// Вариант 5. Выводим Y или P в зависимости от кнопки 0. Кнопка 1 переворачивает букву
// Способ 2. always-блок и оператор 'if'. 
//
//----------------------------------------------------------------------------

module top_5
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    reg [7:1] pio_r;

    always @*
    begin
        if (BTN [1])
        begin
            if (BTN [0])
                pio_r = 7'b0111101;  // перевернутое P
            else
                pio_r = 7'b1010111;  // перевернутое Y
        end
        else
        begin
            if (BTN [0])
                pio_r = 7'b1100111;  // P
            else
                pio_r = 7'b0111011;  // Y
        end
    end
    
    assign pio [7:1] = pio_r;

endmodule

//----------------------------------------------------------------------------
//
// Вариант 6. Выводим Y или P в зависимости от кнопки 0. Кнопка 1 переворачивает букву
// Способ 3. always-блок и оператор 'case'. 
//
//----------------------------------------------------------------------------

module top_6
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    reg [7:1] pio_r;

    always @*
        case (BTN)
        2'b00: pio_r = 7'b0111011;  // Y
        2'b01: pio_r = 7'b1100111;  // P
        2'b10: pio_r = 7'b1010111;  // перевернутое Y
        2'b11: pio_r = 7'b0111101;  // перевернутое P
        endcase
    
    assign pio [7:1] = pio_r;

endmodule

//----------------------------------------------------------------------------
//
// Вариант 7. Выводим числа от 0 до 7 в зависимости от нажатых трех кнопок
//
//----------------------------------------------------------------------------

module top_7
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);
    
    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 7 6 5 4 3 2 1       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 

    wire extra_button = pio [8];
    
    reg [7:1] pio_r;
    
    always @*
        case ( { BTN, extra_button } )
        3'b000: pio_r = 7'b1111110;  // 0 abcdefg
        3'b001: pio_r = 7'b0110000;  // 1
        3'b010: pio_r = 7'b1101101;  // 2
        3'b011: pio_r = 7'b1111001;  // 3
        3'b100: pio_r = 7'b0110011;  // 4
        3'b101: pio_r = 7'b1011011;  // 5
        3'b110: pio_r = 7'b1011111;  // 6
        3'b111: pio_r = 7'b1110000;  // 7
        endcase
    
    assign pio [7:1] = pio_r;

endmodule
