//----------------------------------------------------------------------------
//
//  Пример 1: Простая комбинаторная логика
//
//----------------------------------------------------------------------------

module top
(
    output [1:0] LED,  // Два светодиода
    input  [1:0] BTN   // Две кнопки
);

    assign LED [0] = BTN [0] & BTN [1];
    assign LED [1] = BTN [0] | BTN [1];
    
endmodule
