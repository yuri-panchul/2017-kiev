//----------------------------------------------------------------------------
//
//  Упражнение 14: Мультиплексоры и модули
//
//----------------------------------------------------------------------------

// Выбор одного из двух двухбитовых элементов

module mux_2_1
(
    input  [1:0] d0,
    input  [1:0] d1,
    input        sel,
    output [1:0] y
);

    assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------

// Мультиплексор, выбирающий один из четырех двухбитовых элементов
// Реализация 1 с использованием условного оператора

module mux_4_1_implementation_1
(
    input  [1:0] d0, d1, d2, d3,
    input  [1:0] sel,
    output [1:0] y
);

    assign y = sel [1]
        ? (sel [0] ? d3 : d2)
        : (sel [0] ? d1 : d0);

endmodule

//----------------------------------------------------------------------------

// Мультиплексор, выбирающий один из четырех двухбитовых элементов
// Реализация 2 с использованием оператора выбора case

module mux_4_1_implementation_2
(
    input      [1:0] d0, d1, d2, d3,
    input      [1:0] sel,
    output reg [1:0] y
);

    always @*
        case (sel)
        2'b00: y = d0;
        2'b01: y = d1;
        2'b10: y = d2;
        2'b11: y = d3;
        endcase

endmodule

//----------------------------------------------------------------------------

// Мультиплексор, выбирающий один из четырех двухбитовых элементов
// Реализация 3 с помощью дерева из трех подмодулей с двумя двухбитовыми входами

module mux_4_1_implementation_3
(
    input  [1:0] d0, d1, d2, d3,
    input  [1:0] sel,
    output [1:0] y
);

    wire [1:0] w01, w23;

    mux_2_1 i0 (.d0 ( d0  ), .d1 ( d1  ), .sel (sel [0]), .y ( w01 ));
    mux_2_1 i1 (.d0 ( d2  ), .d1 ( d3  ), .sel (sel [0]), .y ( w23 ));
    mux_2_1 i2 (.d0 ( w01 ), .d1 ( w23 ), .sel (sel [1]), .y ( y   ));

endmodule

//----------------------------------------------------------------------------

// Мультиплексор, выбирающий один из четырех однобитовых элементов

module mux_4_1_bits_1
(
    input        d0, d1, d2, d3,
    input  [1:0] sel,
    output       y
);

    assign y = sel [1]
        ? (sel [0] ? d3 : d2)
        : (sel [0] ? d1 : d0);

endmodule

//----------------------------------------------------------------------------

// Мультиплексор, выбирающий один из четырех двухбитовых элементов
// Реализация 4 с помощью двух подмодулей с четырьмя однобитовыми входами

module mux_4_1_implementation_4
(
    input  [1:0] d0, d1, d2, d3,
    input  [1:0] sel,
    output [1:0] y
);

    mux_4_1_bits_1 high
    (
        .d0  ( d0 [1] ),
        .d1  ( d1 [1] ),
        .d2  ( d2 [1] ),
        .d3  ( d3 [1] ),
        .sel ( sel    ),
        .y   ( y  [1] )
    );

    mux_4_1_bits_1 low
    (
        .d0  ( d0 [0] ),
        .d1  ( d1 [0] ),
        .d2  ( d2 [0] ),
        .d3  ( d3 [0] ),
        .sel ( sel    ),
        .y   ( y  [0] )
    );

endmodule

//----------------------------------------------------------------------------

// Верхний модуль, который устанавливает четыре варианта реализации мультиплексора

module cmod_a7_12
(
    inout  [48:1] pio,  // GPIO, General-Purpose Input/Output
    input  [ 1:0] BTN,  // Две кнопки
    output [ 1:0] LED   // Два светодиода
);

    wire [1:0] d0 = pio [12:11];
    wire [1:0] d1 = pio [14:13];
    wire [1:0] d2 = pio [18:17];
    wire [1:0] d3 = pio [20:19];

    wire [1:0] y0, y1, y2, y3;

    assign pio [8:1] = { y3, y2, y1, y0 };

    assign LED = y0;

    mux_4_1_implementation_1 mux_4_1_i1
    (
        .d0  ( d0  ),
        .d1  ( d1  ),
        .d2  ( d2  ),
        .d3  ( d3  ),
        .sel ( BTN ),
        .y   ( y0  )
    ); 

    mux_4_1_implementation_2 i1
    (
        .d0  ( d0  ),
        .d1  ( d1  ),
        .d2  ( d2  ),
        .d3  ( d3  ),
        .sel ( BTN ),
        .y   ( y1  )
    ); 

    mux_4_1_implementation_3
    (
        .d0  ( d0  ),
        .d1  ( d1  ),
        .d2  ( d2  ),
        .d3  ( d3  ),
        .sel ( BTN ),
        .y   ( y2  )
    ); 

    mux_4_1_implementation_4
    (
        .d0  ( d0  ),
        .d1  ( d1  ),
        .d2  ( d2  ),
        .d3  ( d3  ),
        .sel ( BTN ),
        .y   ( y3  )
    );

endmodule
