//----------------------------------------------------------------------------
//
//  Пример 3: Буква в зависимости от кнопки
//
//----------------------------------------------------------------------------

module top
(
    input  [ 1:0] BTN,         // Две кнопки
    inout  [48:1] pio          // GPIO, General-Purpose Input/Output
);

    // a b c d e f g  dp   Буквы с картинки
    // 7 6 4 2 1 9 10 5    Выводы 7-сегментного индикатора
    // 5 4 3 2 1 6 7       Выводы сигнала pio в ПЛИС
    
    //   --a--
    //  |     |
    //  f     b
    //  |     |
    //   --g--
    //  |     |
    //  e     c
    //  |     |
    //   --d-- 


    // 1. Выводим одну букву Y. Присваиваем по битам.

    /*
    assign pio [1] = 1'b0;  // e
    assign pio [2] = 1'b1;  // d
    assign pio [3] = 1'b1;  // c
    assign pio [4] = 1'b1;  // b
    assign pio [5] = 1'b0;  // a
    assign pio [6] = 1'b1;  // f
    assign pio [7] = 1'b1;  // g
    */
    
    // 2. Выводим одну букву P. Присваиваем целым битовым вектором.

    /*
    assign pio [7:1] = 7'b1111001;  // gfabcde
    */

    // 3. Выводим Y или P в зависимости от кнопки 0.

    `ifdef UNDEF    
    assign pio [7:1] = BTN [0] ? 7'b1111001 /* P */ : 7'b1101110 /* Y */ ;
    `endif

    // 4. Выводим Y или P в зависимости от кнопки 0. Кнопка 1 переворачивает букву

    assign pio [7:1]
        = 
        BTN [1] 
            ? (BTN [0]
                ? 7'b1001111 /* перевернутое P */
                : 7'b1110101 /* перевернутое Y */ )
            : (BTN [0]
                ? 7'b1111001 /* P */
                : 7'b1101110 /* Y */ );

endmodule
