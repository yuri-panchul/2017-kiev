//----------------------------------------------------------------------------
//
//  Пример 1: Простая комбинаторная логика
//
//----------------------------------------------------------------------------

module top
(
    output [1:0] LED,         // Два светодиода

    output       RGB0_Red,    // Красная часть трехцветного светодиода
    output       RGB0_Green,  // Зеленая часть трехцветного светодиода
    output       RGB0_Blue,   // Синяя часть трехцветного светодиода

    input  [1:0] BTN          // Две кнопки
);

    assign LED [0] = BTN [0] & BTN [1];
    assign LED [1] = BTN [0] | BTN [1];

    assign RGB0_Red   = BTN [0];
    assign RGB0_Green = BTN [1];
    assign RGB0_Blue  = BTN [2];
    
endmodule
